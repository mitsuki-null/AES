module Sbox(
    input   [7:0]       IN,
    output  [7:0]       OUT
);

reg         [7:0]       tmp;

always @ (*) begin
    case(IN) begin
        8'h00: tmp<=



    end
end

endmodule